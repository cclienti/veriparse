module repeat1;

  initial
     repeat(10) begin
        $display("repeat!");
     end

endmodule
