module dimension0;
   input reg [3:0] [7:0] a;
   reg [3:0] [4:1] b [0:1] [2:1];
   integer c;
   integer d [7:0];
endmodule
