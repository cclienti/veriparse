/* Module 2 */
module module2(input wire              reset, clk,
               input wire signed [7:0] in0, in1,
               input wire [7:0]        in2, in3,
               output reg              out);
endmodule
