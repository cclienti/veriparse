module block0();
   reg clk,reset,enable,data;

   initial begin
      begin
         clk = 0;
         reset = 0;
      end
      begin
         enable = 0;
         data = 0;
      end
   end

endmodule
