module realconst3
  (input wire        reset,
   input wire        clk,
   input wire [31:0] in,
   output reg [31:0] out);

   always @(posedge clk) out <= 5_0.1_1E+5_0;

endmodule
