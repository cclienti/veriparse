/* Module 0 */
module module0(reset, clk, in0, in1, out);
   input       reset;
   input       clk;
   input [7:0] in0, in1;
   output      out;

   wire        reset, clk;
   wire [7:0]  in0, in1;
endmodule
