module assignment0(input wire  a, b,
                   output wire s);
   always @(*) s = a & b;
endmodule
