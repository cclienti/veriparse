module deadcode7;
   (* ramstyle = "M144K" *) reg [31:0] mem;
   reg test = 0;

   initial begin
      $display(test);
   end
endmodule
