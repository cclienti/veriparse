module instance2;
   my_module inst [3:0] ();
endmodule

module my_module;
endmodule
