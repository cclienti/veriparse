module initial1();
   reg clk, reset, enable, data;

   initial clk = 0;
   initial reset = 0;
   initial enable = 0;
   initial data = 0;

endmodule
