module instance2;
   my_module2 inst [3:0] ();
endmodule

module my_module2;
endmodule
