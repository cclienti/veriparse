module constant_folding1;
   reg [31:0] invert;

   initial begin
      invert = ~(32'h0);
   end

endmodule
