module deadcode4(output reg out0,
                 output out1);
   reg out1;
   reg out2;
endmodule
