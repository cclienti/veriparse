/* Module 1 */
module module1(reset, clk, in0, in1, out);
   input wire              reset, clk;
   input wire signed [7:0] in0, in1;
   output reg              out;
endmodule
