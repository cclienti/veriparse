module var3;

   initial begin
      integer x = 0;
   end

endmodule
