module repeat0;

  initial begin
     repeat(10) begin
        $display("repeat!");
     end
  end

endmodule
